LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.NUMERIC_STD.ALL;

ENTITY MESSAGE_REG_TB IS END ENTITY;

ARCHITECTURE ARCH_MESSAGE_REG_TB OF MESSAGE_REG_TB IS
	COMPONENT MESSAGE_REG IS PORT
	(
		CLK	:IN STD_LOGIC;
		INIT	:IN STD_LOGIC;
		WR		:IN STD_LOGIC;
		ADDR	:IN STD_LOGIC_VECTOR(31 downto 0);
		DIN	:IN STD_LOGIC_VECTOR(31 downto 0);
		DOUT	:OUT STD_LOGIC_VECTOR(127 downto 0)
	);
	END COMPONENT;

	SIGNAL CLK	: STD_LOGIC := '0';
	SIGNAL INIT	: STD_LOGIC := '0';
	SIGNAL WR		: STD_LOGIC := '0';
	SIGNAL ADDR	: STD_LOGIC_VECTOR(31 downto 0) := (OTHERS => '0');
	SIGNAL DIN	: STD_LOGIC_VECTOR(31 downto 0) := (OTHERS => '0');
	SIGNAL DOUT	: STD_LOGIC_VECTOR(127 downto 0) := (OTHERS => '0');
	
	SIGNAL CLKp :time := 40 ns;
BEGIN
	tb: MESSAGE_REG PORT MAP (CLK, INIT, WR, ADDR, DIN, DOUT);

	PROCESS
	BEGIN
		CLK <= '0'; wait for CLKp / 2;
		CLK <= '1'; wait for CLKp / 2;
	END PROCESS;

	PROCESS
	BEGIN
		INIT <= '1'; WR <= '0'; ADDR <= X"00000000"; DIN <= X"00000000"; wait for CLKp;
		INIT <= '0'; WR <= '1'; ADDR <= X"00000004"; DIN <= X"F0000000"; wait for CLKp;
		INIT <= '0'; WR <= '1'; ADDR <= X"00000005"; DIN <= X"0F000000"; wait for CLKp;
		INIT <= '0'; WR <= '1'; ADDR <= X"00000006"; DIN <= X"00F00000"; wait for CLKp;
		INIT <= '0'; WR <= '1'; ADDR <= X"00000007"; DIN <= X"000F0000"; wait for CLKp;

		wait;
	END PROCESS;
END ARCHITECTURE;