LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.STD_LOGIC_UNSIGNED.ALL;
	USE IEEE.NUMERIC_STD.ALL;

ENTITY CONTROL IS
	PORT (
		CLK			:IN STD_LOGIC;
		INIT			:IN STD_LOGIC;
		WR				:IN STD_LOGIC;
		ADDR			:IN STD_LOGIC_VECTOR(31 downto 0);
		DATA_WR		:OUT STD_LOGIC;
		RUN			:OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE ARCH_CONTROL OF CONTROL IS
	SIGNAL COUNTER		:STD_LOGIC_VECTOR(7 downto 0);
BEGIN
	PROCESS(CLK, INIT)
	BEGIN
		IF INIT = '1' THEN
			COUNTER	<= (OTHERS => '0');
		ELSIF CLK = '1' AND CLK'EVENT THEN
			IF (WR = '1' AND ADDR = X"7") OR COUNTER /= X"0" THEN
				IF COUNTER /= X"2C" THEN
					COUNTER	<= COUNTER + 1;
				END IF;
				IF COUNTER = X"2C" THEN
					COUNTER	<= X"00";
				END IF;
			END IF;
		END IF;
	END PROCESS;
	
	RUN		<= '1'
					WHEN COUNTER /= X"0" AND COUNTER /= X"2C"
					ELSE '0';
	DATA_WR	<= '1'
					WHEN COUNTER = X"2C"
					ELSE '0';
END ARCHITECTURE;