LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY KEY_REG IS
	PORT
	(
		CLK	:IN STD_LOGIC;
		INIT	:IN STD_LOGIC;
		WR		:IN STD_LOGIC;
		ADDR	:IN STD_LOGIC_VECTOR(31 downto 0);
		DIN	:IN STD_LOGIC_VECTOR(31 downto 0);
		DOUT	:OUT STD_LOGIC_VECTOR(127 downto 0)
	);
END ENTITY;

ARCHITECTURE ARCH_KEY_REG OF KEY_REG IS
	TYPE MEMORY_BLOCK IS ARRAY (0 to 3) OF STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL KEY		:MEMORY_BLOCK := (OTHERS => (OTHERS => '0'));
BEGIN
	PROCESS(CLK, INIT, KEY)
	BEGIN
		IF INIT = '1' THEN
			KEY	<= (OTHERS => (OTHERS => '0'));
		ELSIF CLK = '1' AND CLK'EVENT THEN
			IF WR = '1' AND ADDR <= X"3" THEN
				KEY(conv_integer(ADDR))	<= DIN;
			END IF;
		END IF;
		
		DOUT	<= KEY(0) & KEY(1) & KEY(2) & KEY(3);
	END PROCESS;
END ARCHITECTURE;