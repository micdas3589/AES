LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY MESSAGE_REG IS
	PORT
	(
		CLK	:IN STD_LOGIC;
		INIT	:IN STD_LOGIC;
		WR		:IN STD_LOGIC;
		ADDR	:IN STD_LOGIC_VECTOR(31 downto 0);
		DIN	:IN STD_LOGIC_VECTOR(31 downto 0);
		DOUT	:OUT STD_LOGIC_VECTOR(127 downto 0)
	);
END ENTITY;

ARCHITECTURE ARCH_MESSAGE_REG OF MESSAGE_REG IS
	TYPE MEMORY_BLOCK IS ARRAY (0 to 3) OF STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL MSG		:MEMORY_BLOCK := (OTHERS => (OTHERS => '0'));
BEGIN
	PROCESS(CLK, INIT, MSG)
	BEGIN
		IF INIT = '1' THEN
			MSG	<= (OTHERS => (OTHERS => '0'));
		ELSIF CLK = '1' AND CLK'EVENT THEN
			IF WR = '1' AND ADDR >= X"4" AND ADDR <= X"7" THEN
				MSG(conv_integer(ADDR)-4)	<= DIN;
			END IF;
		END IF;
		
		DOUT	<= MSG(0) & MSG(1) & MSG(2) & MSG(3);
	END PROCESS;
END ARCHITECTURE;