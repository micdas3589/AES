LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.NUMERIC_STD.ALL;

ENTITY ROUND_TB IS END ENTITY;

ARCHITECTURE ARCH_ROUND_TB OF ROUND_TB IS
	COMPONENT ROUND IS PORT
	(
		CLK			:IN STD_LOGIC;
		INIT			:IN STD_LOGIC;
		RUN_ROUND	:IN STD_LOGIC;
		ROUND_NR		:IN STD_LOGIC_VECTOR(3 downto 0);
		STATE_IN		:IN STD_LOGIC_VECTOR(127 downto 0);
		ROUND_KEY	:IN STD_LOGIC_VECTOR(127 downto 0);
		STATE_OUT	:OUT STD_LOGIC_VECTOR(127 downto 0)
	);
	END COMPONENT;

	SIGNAL CLK			: STD_LOGIC := '0';
	SIGNAL INIT			: STD_LOGIC := '0';
	SIGNAL RUN_ROUND	: STD_LOGIC := '0';
	SIGNAL ROUND_NR		: STD_LOGIC_VECTOR(3 downto 0) := (OTHERS => '0');
	SIGNAL STATE_IN		: STD_LOGIC_VECTOR(127 downto 0) := (OTHERS => '0');
	SIGNAL ROUND_KEY	: STD_LOGIC_VECTOR(127 downto 0) := (OTHERS => '0');
	SIGNAL STATE_OUT	: STD_LOGIC_VECTOR(127 downto 0) := (OTHERS => '0');
	
	SIGNAL CLKp :time := 40 ns;
BEGIN
	tb: ROUND PORT MAP (CLK, INIT, RUN_ROUND, ROUND_NR, STATE_IN, ROUND_KEY, STATE_OUT);

	PROCESS
	BEGIN
		CLK <= '0'; wait for CLKp / 2;
		CLK <= '1'; wait for CLKp / 2;
	END PROCESS;

	PROCESS
	BEGIN
		INIT <= '1'; RUN_ROUND <= '0'; ROUND_NR <= X"0"; STATE_IN <= X"00112233445566778899aabbccddeeff"; ROUND_KEY <= X"000102030405060708090a0b0c0d0e0f"; wait for CLKp;
		INIT <= '0'; RUN_ROUND <= '0'; ROUND_NR <= X"0"; STATE_IN <= X"00112233445566778899aabbccddeeff"; ROUND_KEY <= X"000102030405060708090a0b0c0d0e0f"; wait for CLKp;
		INIT <= '0'; RUN_ROUND <= '1'; ROUND_NR <= X"1"; STATE_IN <= X"00102030405060708090a0b0c0d0e0f0"; ROUND_KEY <= X"d6aa74fdd2af72fadaa678f1d6ab76fe"; wait for 8*CLKp;
		INIT <= '1'; RUN_ROUND <= '0'; ROUND_NR <= X"0"; STATE_IN <= X"00000000000000000000000000000000"; ROUND_KEY <= X"00000000000000000000000000000000"; wait for CLKp;
		INIT <= '0'; RUN_ROUND <= '1'; ROUND_NR <= X"2"; STATE_IN <= X"89d810e8855ace682d1843d8cb128fe4"; ROUND_KEY <= X"b692cf0b643dbdf1be9bc5006830b3fe"; wait for 8*CLKp;
		INIT <= '1'; RUN_ROUND <= '0'; ROUND_NR <= X"0"; STATE_IN <= X"00000000000000000000000000000000"; ROUND_KEY <= X"00000000000000000000000000000000"; wait for CLKp;
		INIT <= '0'; RUN_ROUND <= '1'; ROUND_NR <= X"3"; STATE_IN <= X"4915598f55e5d7a0daca94fa1f0a63f7"; ROUND_KEY <= X"b6ff744ed2c2c9bf6c590cbf0469bf41"; wait for 8*CLKp;
		INIT <= '1'; RUN_ROUND <= '0'; ROUND_NR <= X"0"; STATE_IN <= X"00000000000000000000000000000000"; ROUND_KEY <= X"00000000000000000000000000000000"; wait for CLKp;
		INIT <= '0'; RUN_ROUND <= '1'; ROUND_NR <= X"4"; STATE_IN <= X"fa636a2825b339c940668a3157244d17"; ROUND_KEY <= X"47f7f7bc95353e03f96c32bcfd058dfd"; wait for 8*CLKp;
		INIT <= '1'; RUN_ROUND <= '0'; ROUND_NR <= X"0"; STATE_IN <= X"00000000000000000000000000000000"; ROUND_KEY <= X"00000000000000000000000000000000"; wait for CLKp;
		INIT <= '0'; RUN_ROUND <= '1'; ROUND_NR <= X"5"; STATE_IN <= X"247240236966b3fa6ed2753288425b6c"; ROUND_KEY <= X"3caaa3e8a99f9deb50f3af57adf622aa"; wait for 8*CLKp;
		INIT <= '1'; RUN_ROUND <= '0'; ROUND_NR <= X"0"; STATE_IN <= X"00000000000000000000000000000000"; ROUND_KEY <= X"00000000000000000000000000000000"; wait for CLKp;
		INIT <= '0'; RUN_ROUND <= '1'; ROUND_NR <= X"6"; STATE_IN <= X"c81677bc9b7ac93b25027992b0261996"; ROUND_KEY <= X"5e390f7df7a69296a7553dc10aa31f6b"; wait for 8*CLKp;
		INIT <= '1'; RUN_ROUND <= '0'; ROUND_NR <= X"0"; STATE_IN <= X"00000000000000000000000000000000"; ROUND_KEY <= X"00000000000000000000000000000000"; wait for CLKp;
		INIT <= '0'; RUN_ROUND <= '1'; ROUND_NR <= X"7"; STATE_IN <= X"c62fe109f75eedc3cc79395d84f9cf5d"; ROUND_KEY <= X"14f9701ae35fe28c440adf4d4ea9c026"; wait for 8*CLKp;
		INIT <= '1'; RUN_ROUND <= '0'; ROUND_NR <= X"0"; STATE_IN <= X"00000000000000000000000000000000"; ROUND_KEY <= X"00000000000000000000000000000000"; wait for CLKp;
		INIT <= '0'; RUN_ROUND <= '1'; ROUND_NR <= X"8"; STATE_IN <= X"d1876c0f79c4300ab45594add66ff41f"; ROUND_KEY <= X"47438735a41c65b9e016baf4aebf7ad2"; wait for 8*CLKp;
		INIT <= '1'; RUN_ROUND <= '0'; ROUND_NR <= X"0"; STATE_IN <= X"00000000000000000000000000000000"; ROUND_KEY <= X"00000000000000000000000000000000"; wait for CLKp;
		INIT <= '0'; RUN_ROUND <= '1'; ROUND_NR <= X"9"; STATE_IN <= X"fde3bad205e5d0d73547964ef1fe37f1"; ROUND_KEY <= X"549932d1f08557681093ed9cbe2c974e"; wait for 8*CLKp;
		INIT <= '1'; RUN_ROUND <= '0'; ROUND_NR <= X"0"; STATE_IN <= X"00000000000000000000000000000000"; ROUND_KEY <= X"00000000000000000000000000000000"; wait for CLKp;
		INIT <= '0'; RUN_ROUND <= '1'; ROUND_NR <= X"A"; STATE_IN <= X"bd6e7c3df2b5779e0b61216e8b10b689"; ROUND_KEY <= X"13111d7fe3944a17f307a78b4d2b30c5"; wait for 8*CLKp;
		
		wait;
	END PROCESS;
END ARCHITECTURE;